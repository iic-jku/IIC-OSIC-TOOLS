** sch_path: /foss/pdks/ihp-sg13g2/libs.tech/xschem/sg13g2_tests_xyce/dc_lv_pmos.sch
**.subckt dc_lv_pmos
Vgs GND net1 0
Vds GND net3 0
XM1 net2 net1 GND GND sg13_lv_pmos w=1.0u l=0.45u ng=1
Vd net2 net3 0
**** begin user architecture code
.preprocess replaceground true
.option temp=27
.step  vgs 0.35 1.1 0.05
.dc vds 0 1.2 0.01
.print dc format=raw file=/tmp/dc_lv_pmos.raw i(Vd)
.lib /foss/pdks/ihp-sg13g2/libs.tech/xyce/models/cornerMOSlv.lib mos_tt
**** end user architecture code
**.ends
.GLOBAL GND
.end
